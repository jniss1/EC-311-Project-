`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 12/08/2024 02:45:57 PM
// Design Name: 
// Module Name: memory_module
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module memory_module (
    input wire [9:0] x,         // Current x-coordinate from VGA
    input wire [9:0] y,         // Current y-coordinate from VGA
    output reg [3:0] red,      // 5-bit red color output
    output reg [3:0] green,    // 6-bit green color output
    output reg [3:0] blue      // 5-bit blue color output
);

    // Sprite size
    localparam SPRITE_WIDTH = 64;  // Sprite width (64 pixels)
    localparam SPRITE_HEIGHT = 64; // Sprite height (64 pixels)
    localparam BIT_WIDTH = 12;
    localparam TOTAL_PIXELS = SPRITE_WIDTH * SPRITE_HEIGHT;
    localparam TOTAL_BITS = TOTAL_PIXELS * BIT_WIDTH;

    // Sprite position on the screen
    localparam SPRITE_X_OFFSET = 100; // Horizontal starting position of sprite
    localparam SPRITE_Y_OFFSET = 50;  // Vertical starting position of sprite

    // Memory array for the sprite data
    reg [149151:0] pixel_data;

    // Initialize the memory with data from the .mem file
    initial begin
        pixel_data <= 149151'b000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110111011101001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110111011101010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111110111011101000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100111011101110001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110111111111111100110011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101101110111011110111011101110111011101010001000100000000000000000000000000000000000000000000000000000000000000001100110011000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111111011101110011101110111000100010001000000000000000000000000000000000000000000000000001000100010010101010101101110111011111111111111001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111111011101110010001000100000000000000000000000000000000000000000000000000001000100010101010101010110111011101110111011101100110011001001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001100110011001111011101110010001000100000000000000000000000000000000000000000000000000010101010101111011101110110011001100001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101110111011001100110011011001100110010001000100001000100010011101110111110011001100111011101110011101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100111111111111110011001100110111011101101010101010100010001000111011101110100110011001010001000100000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110111011101011101110111010001000100001100110011000000000000001100110011111011101110100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001001000100010001100110011010001000100011001100110110011001100111111111111001100110011000000000000000000000000000000000000000000000000010101010101111111111111001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001101110111011001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001001000100010001100110011010101010101011101110111100110011001101110111011101110111011110011001100110011001100110011001100110011001100101110111011101010101010100110011001011101110111110011001100011001100110000000000000000000000000000000000000000100010001111011101110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010011101110111011101110111110111011101000100010001000000000000000000000000000000000000000000000000000100010001010001000100011101110111101110111011110111011101110111011101110011001100101110111011100110011001011101110111011001100110010001000100001000100010000100010001000000000000000000000000000000000000000000000000000000000000000000000000011101110111111011101110000100010001000000000000000000000000000000000000100010001000110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011100010001000000000000000101010101010101110111011000100010001010001000100011101110111101110111011110111011101110011001100101010101010011001100110001100110011000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101111111111111000100010001000000000000000000000000000000000000100110011001110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010101110111011000000000000001000100010111011101110111011101110110011001100100110011001011001100110001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010111011101110010101010101000000000000000000000000010101010101111111111111010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001011001100110111011101110001100110011000000000000011001100110111111111111001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110111011101110001000100010000000000000001000100010100010001000101110111011110111011101011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110110011001100110111011101011101110111000000000000000000000000000100010001011101110111110111011101110011001100110111011101011101110111000000000000000000000000110011001100101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101011101110111000000000000000000000000000000000000000000000000010101010101111111111111001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000111011101110010001000100011001100110111011101110001000100010011101110111111011101110110011001100010001000100000000000000010101010101101110111011000000000000000000000000001100110011111011101110001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110111011101100010001000000000000000000000000000000000000000000000000000001000100010111011101110010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001111011101110011001100110000000000000001000100010111111111111111011101110110011001100010101010101000000000000000000000000000000000000000100010001110011001100001000100010000000000000000000000000100110011001101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001010001000100000000000000000000000000000000000000000000000000010101010101111011101110000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110111011101010101010101000000000000100110011001111011101110011101110111000000000000000000000000000000000000000000000000000000000000000000000000101010101010010001000100000000000000000000000000010001000100111111111111010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101010101010101000000000000000000000000000000000000001100110011111011101110001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111111011101110110111011101110111011101001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110100110011001011001100110110011001100111111111111111111111111110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010011001100110000000000000000000000000000000000000110111011101011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100111111111111101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010111111111111111111111111111111111111110011001100100010001000111111111111010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001001100110011010001000100001100110011010101010101111011101110001000100010000000000000000000000000110011001100011101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101111111111111011101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100100110011001001100110011000000000000000000000000100110011001110111011101000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010100110011001110111011101111111111111111111111111111111111111111111111111111111111111100110011001000000000000000000000000110011001100011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011111111111111011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001011001100110000000000000000000000000000000000000001000100010111111111111011101110111000000000000000000000000000000000000000000000000000000000000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101000000000000000000000000110011001100011101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100101110111011000000000000000000000000000000000000000000000000101110111011111011101110000100010001000000000000000000000000010101010101101110111011111011101110010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110011001100001100110011000000000000000000000000110111011101011001100110000000000000000000000000000000000000000000000000000000000000000000000000001100110011010101010101011101110111101010101010000000000000010001000100111111111111001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011001100110011000000000000000000000000011001100110111111111111111011101110001000100010000000000000100110011001111111111111111111111111111111111111011101110111000000000000000000000000000000000000000000000000000000000000000000000000011001100110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101110111011000100010001000000000000000000000000000100010001111011101110010101010101000000000000010101010101011101110111100010001000100010001000110011001100110011001100100010001000011101110111011001100110000000000000101010101010110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110100110011001000100010001100110011001111111111111110011001100001000100010000000000000011101110111111111111111111111111111111111111111111111111111010001000100000000000000000000000000000000000000000000000000000000000000001000100010111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001000100000000000000000000000000000000000000000100010001101110111011010101010101011101110111011101110111011001100110011101110111101110111011100110011001000000000000000000000000000000000000000000000000000000000000110011001100100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010111011101110111011101110111111111111100010001000000000000000001100110011100010001000010101010101111111111111111111111111111111111111011101110111000000000000000000000000000000000000000000000000000000000000000000000000100010001000111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001100110011000000000000000000000000000000000000000000000000000100010001011001100110100110011001100010001000011101110111100010001000010101010101000000000000000000000000000000000000000000000000000000000000001000100010111111111111010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011111111111111010001000100000000000000000000000000110111011101111011101110001100110011110111011101101110111011010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000110011001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010101010101000000000000000000000000000000000000000000000000011101110111101110111011010101010101001100110011001100110011000100010001000000000000000000000000000000000000000000000000000000000000000000000000010101010101111011101110000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010110111011101111111111111101110111011000100010001001000100010111111111111110011001100000100010001010001000100001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111000000000000000000000000000000000000001000100010000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110110111011101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110111011101101010101010101010101010111111111111110011001100000100010001100110011001011001100110100010001000111111111111111011101110011101110111000000000000000000000000000000000000000000000000000000000000000000000000001100110011111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101010000000000000000000000000000000000000011101110111010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100111011101110000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101110111011000000000000000000000000100010001000111111111111110111011101001100110011010001000100111111111111111111111111111111111111111111111111100010001000000000000000000000000000000000000000000000000000000000000000001000100010111011101110111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110000100010001000000000000000000000000101010101010010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011111111111111001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001101110111011000000000000000000000000000000000000001000100010111011101110111111111111010001000100000100010001111011101110111111111111111111111111111111111111111111111111010001000100000000000000000000000000000000000000000000000000000000000000110111011101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111110111011101000000000000000000000000000100010001110111011101001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001111011101110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010110111011101000100010001000000000000000000000000001000100010110111011101110111011101001100110011000000000000000000000000010101010101111111111111111111111111111111111111111111111111100010001000000000000000000000000000000000000000000000000000000000000000100110011001111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111011101110111000000000000000000000000000000000000101110111011101010101010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101110111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010111011101110001000100010000000000000000000000000010001000100111011101110101110111011000100010001000000000000000000000000000000000000000000000000011001100110111111111111111111111111111111111111110011001100000000000000000000000000000000000000000000000000000000000000010101010101111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111001000100010000000000000000000000000000000000000001000100010111011101110011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011111011101110010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110111111111111010001000100000000000000000000000000011101110111111111111111011101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011110011001100111111111111101010101010000000000000000000000000000000000000000000000000000000000000000100010001110011001100111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111010001000100000000000000000000000000000000000000000000000000011001100110111011101110000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000110111011101000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010111011101110011001100110000000000000000100010001101010101010111011101110010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010000100010001000000000000000000000000000000000000000000000000000000000000000000000000000100010001101010101010111111111111111111111111111111111111111111111111111111111111111111111111111111111111101010101010000000000000000000000000000000000000000000000000000100010001110111011101011101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011100110011001110011001100101110111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011100010001000000000000000001100110011110111011101101110111011000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011100010001000110011001100110111011101110111011101101110111011110011001100111011101110000100010001000000000000000000000000000000000000000000000000100110011001110011001100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010110111011101010001000100000000000000110011001100101110111011000100010001000000000000000000000000000000000000000000000000100110011001100110011001000000000000010101010101111011101110100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001111011101110010001000100000000000000000000000000000000000000000000000000010101010101111011101110000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001000101110111011000000000000000000000000000100010001111011101110111011101110011001100110000000000000000000000000011001100110101010101010000000000000100010001000111011101110010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000111011101110011001100110000000000000000000000000000000000000000100010001010001000100100010001000100110011001101010101010101010101010110011001100110011001100011101110111001000100010000000000000000000000000110011001100100010001000000000000000000000000000011001100110110111011101010101010101110011001100110011001100011101110111011101110111001000100010101110111011110011001100001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011111111111111010001000100000000000000000000000000001100110011101110111011001000100010000000000000000100010001001100110011010001000100001100110011010101010101101110111011011001100110000000000000000000000000100110011001101110111011000000000000000000000000110111011101011001100110000000000000000000000000011001100110110111011101010101010101111011101110101010101010000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110111011101100110011001000000000000000000000000010101010101110111011101010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010110111011101101110111011100010001000111011101110001000100010000000000000000000000000010101010101111111111111100010001000011101110111110011001100110111011101011101110111001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010001000100110111011101101010101010000000000000000000000000001000100010111111111111010101010101000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001011001100110100110011001010101010101000000000000000000000000000000000000000100010001001000100010000000000000000000000000000000000000010001000100101010101010110111011101101010101010010001000100000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010110011001100110111011101011101110111000000000000000000000000001100110011110011001100101110111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001011001100110110011001100110011001100100110011001010001000100000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010110011001100000000000000000000000000000000000000011001100110111011101110100010001000000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011100010001000101110111011110011001100101010101010011101110111010001000100001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001010101010101111011101110010001000100000000000000000000000000011001100110111111111111010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001100110011011001100110100110011001101110111011110011001100101110111011101010101010100010001000010001000100001000100010000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100110011001110111011101101110111011011001100110000000000000000000000000000000000000010001000100111011101110010001000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001010001000100011001100110100010001000101110111011110011001100110011001100110011001100101110111011101010101010100110011001100010001000011001100110100010001000111011101110001000100010000000000000000000000000000000000000000000000000000000000000000000000000110011001100100110011001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001001100110011010001000100010101010101101010101010011101110111100110011001101110111011011101110111000000000000000000000000010001000100011001100110011101110111010101010101011001100110111111111111011001100110000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010101010101011101110111000000000000000000000000000000000000000000000000100110011001110011001100010101010101001100110011000100010001000000000000001100110011100110011001110011001100100010001000011001100110011001100110010101010101001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101010101010101010101010000000000000001000100010100110011001111011101110001000100010000000000000000000000000000000000000000000000000000000000000000000000000001100110011011101110111100110011001101010101010101010101010110111011101101010101010000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011110111011101110011001100100110011001001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000100010100110011001001100110011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001111011101110100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011001100110111011101110000100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001111011101110011101110111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000011101110111111011101110001000100010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000101110111011101110111011000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100010001110011001100100010001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
    end

    // Determine if the current VGA coordinates are within the sprite's bounds
    wire sprite_active = (x >= SPRITE_X_OFFSET && x < SPRITE_X_OFFSET + SPRITE_WIDTH) &&
                         (y >= SPRITE_Y_OFFSET && y < SPRITE_Y_OFFSET + SPRITE_HEIGHT);

    // Calculate pixel index relative to the sprite's top-left corner
    wire [5:0] sprite_x = x - SPRITE_X_OFFSET; // Sprite-relative X coordinate
    wire [5:0] sprite_y = y - SPRITE_Y_OFFSET; // Sprite-relative Y coordinate
    wire [11:0] pixel_index = sprite_y * SPRITE_WIDTH + sprite_x;

    // Output pixel data
    // wire [15:0] pixel_value = sprite_active ? pixel_data[pixel_index] : 16'b0;

   
    
    always @(*)
    begin
        if(sprite_active) begin
            // Extract RGB565 components
            red = pixel_data[(pixel_index*12+8)+:4];
            green = pixel_data[(pixel_index*12+4)+:4]; 
            blue  = pixel_data[(pixel_index*12)+:4];
        end 
        else begin 
            red <= 0;
            green <= 4'b0;
            blue <= 4'b0;
        end
    end

endmodule
